//////////////////////////////////////////////////
// Title:   testPr_hdlc
// Author: 
// Date:  
//////////////////////////////////////////////////

/* testPr_hdlc contains the simulation and immediate assertion code of the
   testbench. 

   For this exercise you will write immediate assertions for the Rx module which
   should verify correct values in some of the Rx registers for:
   - Normal behavior
   - Buffer overflow 
   - Aborts

   HINT:
   - A ReadAddress() task is provided, and addresses are documentet in the 
     HDLC Module Design Description
*/

program testPr_hdlc(
  in_hdlc uin_hdlc
);
  
  int TbErrorCnt;

  // HDLC register addresses:
  const logic [2:0] RX_BUFFER_ADDR = 3'b011;
  const logic [2:0] RXSC = 3'b010;

  /****************************************************************************
   *                                                                          *
   *                               Student code                               *
   *                                                                          *
   ****************************************************************************/

  `include "hdlc_shared.sv"

  // VerifyAbortReceive should verify correct value in the Rx status/control
  // register, and that the Rx data buffer is zero after abort.
  task VerifyAbortReceive(logic [127:0][7:0] data, int Size);
    logic [7:0] ReadData;

    //Verify status register bits
    ReadAddress(Rx_SC, ReadData);
    // INSERT CODE HERE
    assert (ReadData[Rx_Ready] == 1)
      $display("ABORT_RECEIVE: ERROR: Rx_ready should not be high");
    else
      $display("ABORT_RECEIVE:: SUCCESS: Rx_ready is low");

    assert (ReadData[Rx_FrameError] == 1)
      $display("ABORT_RECEIVE: ERROR: Rx_FrameError should not be high");
    else
      $display("ABORT_RECEIVE:: SUCCESS: Rx_FrameError is low");

    assert (ReadData[Rx_Overflow] == 1)
      $display("ABORT_RECEIVE: ERROR: Rx_Overflow should not be high");
    else
      $display("ABORT_RECEIVE:: SUCCESS: Rx_Overflow is low");

    assert (ReadData[Rx_AbortSignal] == 1)
      $display("ABORT_RECEIVE:: SUCCESS: Rx_FrameError is low");
    else
      $display("ABORT_RECEIVE: ERROR: Rx_AbortSignal should not be low");
    
     // Verify all bytes from the Rx_Buff are zero
     for (int i = 0; i < Size; i++) begin
        ReadAddress(RX_BUFFER_ADDR, ReadData);
        assert (ReadData == 0)
            $display("SUCCESS: Rx_Buff is empty: ReadData = %0h", ReadData);
        else
            $display("ERROR: Rx_Buff is not empty: ReadData = %0h", ReadData);
    end

  endtask

  // VerifyNormalReceive should verify correct value in the Rx status/control
  // register, and that the Rx data buffer contains correct data.
  task VerifyNormalReceive(logic [127:0][7:0] data, int Size);
    logic [7:0] ReadData;
    wait(uin_hdlc.Rx_Ready);
    //Verify status register bits
    ReadAddress(Rx_SC, ReadData);

    // INSERT CODE HERE
    assert (ReadData[Rx_Overflow] == 1)
      $display("NORMAL RECEIVE:: ERROR: x OVERFLOW DETECTED!\n");
    else
      $display("NORMAL RECEIVE: SUCCESS: No Rx overflow detected\n");

    assert (ReadData[Rx_AbortSignal] == 1)
      $display("NORMAL RECEIVE:: ERROR: Rx ABORT DETECTED!\n");
    else
      $display("NORMAL RECEIVE:: SUCCESS: No Rx abort detected\n");

    assert (ReadData[Rx_FrameError] == 1)
      $display("NORMAL RECEIVE:: ERROR: INVALID Rx FRAME DETECTED!\n");
    else
      $display("NORMAL RECEIVE:: SUCCESS: FRAME IS VALID\n");

    assert (ReadData[Rx_Ready] == 1)
      $display("NORMAL RECEIVE:: SUCCESS: Rx BUFFER IS READY\n");
    else
      $display("NORMAL RECEIVE:: ERROR: Rx BUFFER NOT READY\n");

    // Verify all bytes from the Rx_Buff
    for (int i = 0; i < Size; i++) begin
        ReadAddress(RX_BUFFER_ADDR, ReadData);
        assert (data[i] == ReadData)
            $display("Rx_Buff has correct data at index %0d: data[%0d] = %0h, ReadData = %0h", 
                      i, i, data[i], ReadData);
        else
            $display("DATA ERROR: Mismatch at index %0d: data[%0d] = %0h, ReadData = %0h", 
                    i, i, data[i], ReadData);
    end
  
  endtask

  // VerifyNormalReceive should verify correct value in the Rx status/control
  // register, and that the Rx data buffer contains correct data.
  task VerifyOverflowReceive(logic [127:0][7:0] data, int Size);
    logic [7:0] ReadData;

     // Verify status register bits
    ReadAddress(Rx_SC, ReadData);

    // INSERT CODE HERE
    assert (ReadData[Rx_Ready] == 1)
      $display("OVERFLOW_RECEIVE:: SUCCESS: Rx_ready is high");
    else
      $display("OVERFLOW_RECEIVE:: ERROR: Rx_ready should not be low");

    assert (ReadData[Rx_FrameError] == 1)
      $display("OVERFLOW_RECEIVE: ERROR: Rx_FrameError should not be high");
    else
      $display("OVERFLOW_RECEIVE:: SUCCESS: Rx_FrameError is low");

    assert (ReadData[Rx_Overflow] == 1)
      $display("OVERFLOW_RECEIVE:: SUCCESS: Rx_Overflow is high");
    else
      $display("OVERFLOW_RECEIVE:: ERROR: Rx_Overflow is low");

    assert (ReadData[Rx_AbortSignal] == 1)
      $display("OVERFLOW_RECEIVE:: ERROR: Rx_AbortSignal should not be low");
    else
      $display("OVERFLOW_RECEIVE: SUCCESS: Rx_AbortSignal is low");
  
  endtask

  //Verify error receive checks all flags correct and Rx_Buff is empty
  task VerifyErrorReceive(logic [127:0][7:0] data, int Size);
    logic [7:0] ReadData;

    // Verify status register bits
    ReadAddress(Rx_SC, ReadData);

    //Might be overkill to check all of these 
    assert (ReadData[Rx_Ready] == 0)
      $display("ERROR_RECEIVE:: SUCCESS: Rx_Ready is low after error");  
    else
      $display("ERROR_RECEIVE:: ERROR: Rx_Ready is high after error");

    assert (ReadData[Rx_FrameError] == 1)
      $display("ERROR_RECEIVE:: SUCCESS: Rx_FrameError is high after error");
    else
      $display("ERROR_RECEIVE:: ERROR: Rx_FrameError is low after error");

    assert (ReadData[Rx_Overflow] == 0)
      $display("ERROR_RECEIVE:: SUCCESS: Rx_Overflow is low after error");
    else
      $display("ERROR_RECEIVE:: ERROR: Rx_Overflow is high after error");

    assert (ReadData[Rx_AbortSignal] == 0)
      $display("ERROR_RECEIVE:: SUCCESS: Rx_AbortSignal is low after error");
    else
      $display("ERROR_RECEIVE:: ERROR: Rx_AbortSignal is high after error");

    assert (ReadData[Rx_Drop] == 0)
      $display("ERROR_RECEIVE:: SUCCESS: Rx_Drop is low after error");
    else
      $display("ERROR_RECEIVE:: ERROR: Rx_Drop is high after error");
    
     // Verify all bytes from the Rx_Buff are zero
     for (int i = 0; i < Size; i++) begin
        ReadAddress(RX_BUFFER_ADDR, ReadData);
        assert (ReadData == 0)
            $display("ERROR_RECEIVE:: SUCCESS: Rx_Buff is empty: ReadData = %0h", ReadData);
        else
            $display("ERROR_RECEIVE:: ERROR: Rx_Buff is not empty: ReadData = %0h", ReadData);
    end
  endtask

  task VerifyDropReceive(logic [127:0][7:0] data, int Size);
    logic [7:0] ReadData;
    // Verify status register bits
    ReadAddress(Rx_SC, ReadData);
    //Check all flags
    assert (ReadData[Rx_Ready] == 0)
      $display("DROP_RECEIVE:: SUCCESS: Rx_Ready is low after dropped frame");
    else
      $display("DROP_RECEIVE:: ERROR: Rx_Ready is high after dropped frame");

    assert (ReadData[Rx_FrameError] == 0)
      $display("DROP_RECEIVE:: SUCCESS: Rx_FrameError is low after dropped frame");
    else
      $display("DROP_RECEIVE:: ERROR: Rx_FrameError is high after dropped frame");

    assert (ReadData[Rx_Overflow] == 0)
      $display("DROP_RECEIVE:: SUCCESS: Rx_Overflow is low after dropped frame");
    else
      $display("DROP_RECEIVE:: ERROR: Rx_Overflow is high after dropped frame");

    assert (ReadData[Rx_AbortSignal] == 0)
      $display("DROP_RECEIVE:: SUCCESS: Rx_AbortSignal is low after dropped frame");
    else
      $display("DROP_RECEIVE:: ERROR: Rx_AbortSignal is high after dropped frame");

    // Verify all bytes from the Rx_Buff are zero
     for (int i = 0; i < Size; i++) begin
        ReadAddress(RX_BUFFER_ADDR, ReadData);
        assert (ReadData == 0)
            $display("DROP_RECEIVE:: SUCCESS: Rx_Buff is empty: ReadData = %0h", ReadData);
        else
            $display("DROP_RECEIVE:: ERROR: Rx_Buff is not empty: ReadData = %0h", ReadData);
    end

  endtask
  
  /****************************************************************************
   *                                                                          *
   *                             Simulation code                              *
   *                                                                          *
   ****************************************************************************/

  initial begin
    $display("*************************************************************");
    $display("%t - Starting Test Program", $time);
    $display("*************************************************************");

    Init();

    //Receive: Size, Abort, FCSerr, NonByteAligned, Overflow, Drop, SkipRead
    Receive( 10, 0, 0, 0, 0, 0, 0); //Normal
    Receive( 40, 1, 0, 0, 0, 0, 0); //Abort
    Receive(126, 0, 0, 0, 1, 0, 0); //Overflow
    Receive( 45, 0, 0, 0, 0, 0, 0); //Normal
    Receive(126, 0, 0, 0, 0, 0, 0); //Normal
    Receive(122, 1, 0, 0, 0, 0, 0); //Abort
    Receive(126, 0, 0, 0, 1, 0, 0); //Overflow
    Receive( 25, 0, 0, 0, 0, 0, 0); //Normal
    Receive( 47, 0, 0, 0, 0, 0, 0); //Normal
    Receive( 42, 0, 0, 0, 0, 1, 0); //FrameDropped
    Receive( 14, 0, 0, 0, 0, 0, 0); //Normal
    Receive( 14, 0, 0, 1, 0, 0, 0); //NonByteAligned
    Receive( 14, 0, 1, 0, 0, 0, 0); //FCSerr

    $display("*************************************************************");
    $display("%t - Finishing Test Program", $time);
    $display("*************************************************************");
    $stop;
  end

  final begin

    $display("*********************************");
    $display("*                               *");
    $display("* \tAssertion Errors: %0d\t  *", TbErrorCnt + uin_hdlc.ErrCntAssertions);
    $display("*                               *");
    $display("*********************************");

  end

  task Init();
    uin_hdlc.Clk         =   1'b0;
    uin_hdlc.Rst         =   1'b0;
    uin_hdlc.Address     = 3'b000;
    uin_hdlc.WriteEnable =   1'b0;
    uin_hdlc.ReadEnable  =   1'b0;
    uin_hdlc.DataIn      =     '0;
    uin_hdlc.TxEN        =   1'b1;
    uin_hdlc.Rx          =   1'b1;
    uin_hdlc.RxEN        =   1'b1;

    TbErrorCnt = 0;

    #1000ns;
    uin_hdlc.Rst         =   1'b1;
  endtask

  task WriteAddress(input logic [2:0] Address ,input logic [7:0] Data);
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Address     = Address;
    uin_hdlc.WriteEnable = 1'b1;
    uin_hdlc.DataIn      = Data;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.WriteEnable = 1'b0;
  endtask

  task ReadAddress(input logic [2:0] Address ,output logic [7:0] Data);
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Address    = Address;
    uin_hdlc.ReadEnable = 1'b1;
    #100ns;
    Data                = uin_hdlc.DataOut;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.ReadEnable = 1'b0;
  endtask

  task InsertFlagOrAbort(int flag);
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b0;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b1;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b1;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b1;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b1;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b1;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b1;
    @(posedge uin_hdlc.Clk);
    if(flag)
      uin_hdlc.Rx = 1'b0;
    else
      uin_hdlc.Rx = 1'b1;
  endtask

  task MakeRxStimulus(logic [127:0][7:0] Data, int Size);
    logic [4:0] PrevData;
    PrevData = '0;
    for (int i = 0; i < Size; i++) begin
      for (int j = 0; j < 8; j++) begin
        if(&PrevData) begin
          @(posedge uin_hdlc.Clk);
          uin_hdlc.Rx = 1'b0;
          PrevData = PrevData >> 1;
          PrevData[4] = 1'b0;
        end

        @(posedge uin_hdlc.Clk);
        uin_hdlc.Rx = Data[i][j];

        PrevData = PrevData >> 1;
        PrevData[4] = Data[i][j];
      end
    end
  endtask

  task Receive(int Size, int Abort, int FCSerr, int NonByteAligned, int Overflow, int Drop, int SkipRead);
    logic [127:0][7:0] ReceiveData;
    logic       [15:0] FCSBytes;
    logic   [2:0][7:0] OverflowData;
    string msg;
    if(Abort)
      msg = "- Abort";
    else if(FCSerr)
      msg = "- FCS error";
    else if(NonByteAligned)
      msg = "- Non-byte aligned";
    else if(Overflow)
      msg = "- Overflow";
    else if(Drop)
      msg = "- Drop";
    else if(SkipRead)
      msg = "- Skip read";
    else
      msg = "- Normal";
    $display("*************************************************************");
    $display("%t - Starting task Receive %s", $time, msg);
    $display("*************************************************************");

    for (int i = 0; i < Size; i++) begin
      ReceiveData[i] = $urandom;
    end
    ReceiveData[Size]   = '0;
    ReceiveData[Size+1] = '0;

    //Calculate FCS bits;
    GenerateFCSBytes(ReceiveData, Size, FCSBytes);
    ReceiveData[Size]   = FCSBytes[7:0];
    ReceiveData[Size+1] = FCSBytes[15:8];

    //Enable FCS
    if(!Overflow && !NonByteAligned)
      WriteAddress(RXSC, 8'h20);
    else
      WriteAddress(RXSC, 8'h00);

     if(FCSerr) begin
      ReceiveData[Size-1] -= 1;
    end


    //Generate stimulus
    InsertFlagOrAbort(1);
    
    MakeRxStimulus(ReceiveData, Size + 2);
    
    if(Overflow) begin
      OverflowData[0] = 8'h44;
      OverflowData[1] = 8'hBB;
      OverflowData[2] = 8'hCC;
      MakeRxStimulus(OverflowData, 3);
    end

    if (NonByteAligned) begin
      @(posedge uin_hdlc.Clk);
      uin_hdlc.Rx = 0;
    end

    if(Abort) begin
      InsertFlagOrAbort(0);
    end else begin
      InsertFlagOrAbort(1);
    end

    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b1;

    repeat(8)
      @(posedge uin_hdlc.Clk);

    if(Drop) begin 
      WriteAddress(Rx_SC, 8'b1 << Rx_Drop);
    end
    
    if(Abort)
      VerifyAbortReceive(ReceiveData, Size);
    else if(Overflow)
      VerifyOverflowReceive(ReceiveData, Size);
    else if(Drop)
      VerifyDropReceive(ReceiveData, Size);
    else if(FCSerr || NonByteAligned)
      VerifyErrorReceive(ReceiveData, Size);
    else if(!SkipRead)
      VerifyNormalReceive(ReceiveData, Size);

    #5000ns;
  endtask

  task GenerateFCSBytes(logic [127:0][7:0] data, int size, output logic[15:0] FCSBytes);
    logic [23:0] CheckReg;
    CheckReg[15:8]  = data[1];
    CheckReg[7:0]   = data[0];
    for(int i = 2; i < size+2; i++) begin
      CheckReg[23:16] = data[i];
      for(int j = 0; j < 8; j++) begin
        if(CheckReg[0]) begin
          CheckReg[0]    = CheckReg[0] ^ 1;
          CheckReg[1]    = CheckReg[1] ^ 1;
          CheckReg[13:2] = CheckReg[13:2];
          CheckReg[14]   = CheckReg[14] ^ 1;
          CheckReg[15]   = CheckReg[15];
          CheckReg[16]   = CheckReg[16] ^1;
        end
        CheckReg = CheckReg >> 1;
      end
    end
    FCSBytes = CheckReg;
  endtask

endprogram
